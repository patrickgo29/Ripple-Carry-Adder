library verilog;
use verilog.vl_types.all;
entity fourbitRCAdder_vlg_vec_tst is
end fourbitRCAdder_vlg_vec_tst;
